-- pong.vhdl
-- Tarrin Rasmussen 11/18/2019