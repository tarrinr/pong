pll_adc_inst : pll_adc PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		locked	 => locked_sig
	);
